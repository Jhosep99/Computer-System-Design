library verilog;
use verilog.vl_types.all;
entity Outs_16_Ports_vlg_vec_tst is
end Outs_16_Ports_vlg_vec_tst;
